--+----------------------------------------------------------------------------
--| 
--| DESCRIPTION   : This file implements the top level module for a BASYS 
--|
--|     Ripple-Carry Adder: S = A + B
--|
--|     Our **user** will input the following:
--|
--|     - $C_{in}$ on switch 0
--|     - $A$ on switches 4-1
--|     - $B$ on switches 15-12
--|
--|     Our **user** will expect the following outputs:
--|
--|     - $Sum$ on LED 3-0
--|     - $C_{out} on LED 15
--|
--+----------------------------------------------------------------------------
--|
--| NAMING CONVENSIONS :
--|
--|    xb_<port name>           = off-chip bidirectional port ( _pads file )
--|    xi_<port name>           = off-chip input port         ( _pads file )
--|    xo_<port name>           = off-chip output port        ( _pads file )
--|    b_<port name>            = on-chip bidirectional port
--|    i_<port name>            = on-chip input port
--|    o_<port name>            = on-chip output port
--|    c_<signal name>          = combinatorial signal
--|    f_<signal name>          = synchronous signal
--|    ff_<signal name>         = pipeline stage (ff_, fff_, etc.)
--|    <signal name>_n          = active low signal
--|    w_<signal name>          = top level wiring signal
--|    g_<generic name>         = generic
--|    k_<constant name>        = constant
--|    v_<variable name>        = variable
--|    sm_<state machine type>  = state machine type definition
--|    s_<signal name>          = state name
--|
--+----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;


entity top_basys3 is
	port(
		-- Switches
		sw		:	in  std_logic_vector(15 downto 0);
		
		-- LEDs
		led	    :	out	std_logic_vector(15 downto 0)
	);
end top_basys3;

architecture top_basys3_arch of top_basys3 is 
	component ripple_adder is
    Port ( A : in STD_LOGIC_VECTOR (3 downto 0);
           B : in STD_LOGIC_VECTOR (3 downto 0);
           Cin : in STD_LOGIC;
           S : out STD_LOGIC_VECTOR (3 downto 0);
           Cout : out STD_LOGIC);
    end component;
    -- declare the component of your top-level design

    -- declare any signals you will need
    signal w_sw0 : std_logic := '0';
    signal w_sw1 : std_logic := '0';
    signal w_sw2 : std_logic := '0';
    signal w_sw3 : std_logic := '0';
    signal w_sw4 : std_logic := '0';
    signal w_sw12 : std_logic := '0';
    signal w_sw13 : std_logic := '0';
    signal w_sw14 : std_logic := '0';
    signal w_sw15 : std_logic := '0';
    signal w_led0 : std_logic := '0';
    signal w_led1 : std_logic := '0';
    signal w_led2 : std_logic := '0';
    signal w_led3 : std_logic := '0';
    signal w_led15 : std_logic := '0';
  
begin
	-- PORT MAPS --------------------
   ripple_inst : ripple_adder port map(
    A(0) => w_sw1,
    A(1) => w_sw2,
    A(2) => w_sw3,
    A(3) => w_sw4,
    B(0) => w_sw12,
    B(1) => w_sw13,
    B(2) => w_sw14,
    B(3) => w_sw15,
    Cin  => w_sw0,
    S(0) => w_led0,
    S(1) => w_led1,
    S(2) => w_led2,
    S(3) => w_led3,
    Cout => w_led15
   );
	---------------------------------
	
	-- CONCURRENT STATEMENTS --------
	led(14 downto 4) <= (others => '0'); -- Ground unused LEDs
	w_sw0  <= sw(0);
    w_sw1  <= sw(1);
    w_sw2  <= sw(2);
    w_sw3  <= sw(3);
    w_sw4  <= sw(4);
    w_sw12 <= sw(12);
    w_sw13 <= sw(13);
    w_sw14 <= sw(14);
    w_sw15 <= sw(15);
    led(0)  <= w_led0;
    led(1)  <= w_led1;
    led(2)  <= w_led2;
    led(3)  <= w_led3;
    led(15) <= w_led15;
	---------------------------------
end top_basys3_arch;
